module xor_gate();
initial
$display("hello");
endmodule

